//
// Copyright (C) 2008 Intel Corporation
//
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
//

// Simulation Physical Platform

import Clocks::*;
import Vector::*;

`include "clocks_device.bsh"
`include "unix_comm_device.bsh"
`include "physical_platform_utils.bsh"

// PHYSICAL_DRIVERS

// This represents the collection of all platform capabilities which the
// rest of the FPGA uses to interact with the outside world.
// We use other modules to actually do the work.

interface PHYSICAL_DRIVERS;

    interface CLOCKS_DRIVER    clocksDriver;
    interface Vector#(`NUM_FPGA,UNIX_COMM_DRIVER) unixCommDrivers;

endinterface

// TOP_LEVEL_WIRES

// The TOP_LEVEL_WIRES is the datatype which gets passed to the top level
// and output as input/output wires. These wires are then connected to
// physical pins on the FPGA as specified in the accompanying UCF file.
// These wires are defined in the individual devices.

interface TOP_LEVEL_WIRES;
    
    interface CLOCKS_WIRES    clocksWires;
    interface Vector#(`NUM_FPGA, UNIX_COMM_WIRES) unixCommWires;
    
endinterface

// PHYSICAL_PLATFORM

// The platform is the aggregation of wires and drivers.

interface PHYSICAL_PLATFORM;
    
    interface PHYSICAL_DRIVERS physicalDrivers;
    interface TOP_LEVEL_WIRES  topLevelWires;

endinterface

// mkPhysicalPlatform

// This is a convenient way for the outside world to instantiate all the devices
// and an aggregation of all the wires.

module mkPhysicalPlatform
    // interface:
    (PHYSICAL_PLATFORM);
    
    // The Platform is instantiated inside a NULL clock domain. Our first course of
    // action should be to instantiate the Clocks Physical Device and obtain interfaces
    // to clock and reset the other devices with.
    
    CLOCKS_DEVICE clocks_device <- mkClocksDevice();
    
    Clock clk = clocks_device.driver.clock;
    Reset rst = clocks_device.driver.reset;
    
    Vector#(`NUM_FPGA, UNIX_COMM_DRIVER) unixDrivers = newVector();
    Vector#(`NUM_FPGA, UNIX_COMM_WIRES)  unixWires = newVector();
    for(Integer i = 0; i < `NUM_FPGA; i = i +1)
    begin 
        if(i != `MY_ID)
        begin
	   let dev <- mkUNIXCommDevice("/tmp/FPGA" + integerToString(`MY_ID) +"ToFPGA" + integerToString(i),
                                       "/tmp/FPGA" + integerToString(i) + "ToFPGA" + integerToString(`MY_ID),
                                       clocked_by clk,
                                       reset_by rst);
           unixDrivers[i] = dev.driver;
           unixWires[i]   = dev.wires;
        end
    end 

    // Finally, instantiate all other physical devices

    // Aggregate the drivers
    
    interface PHYSICAL_DRIVERS physicalDrivers;
    
        interface clocksDriver   = clocks_device.driver;
        interface unixCommDrivers = unixDrivers;

    endinterface
    
    // Aggregate the wires
    
    interface TOP_LEVEL_WIRES topLevelWires;
    
        interface clocksWires    = clocks_device.wires;
        interface unixCommWires  = unixWires;

    endinterface
               
endmodule
