`include "asim/provides/soft_connections.bsh"
`include "asim/provides/test_d.bsh"

module [CONNECTED_MODULE] mkB (Empty);
    let d <- mkD();
endmodule

