//
// Copyright (C) 2008 Intel Corporation
//
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
//

import FIFOF::*;
import Vector::*;
import GetPut::*;
import Connectable::*;
import Clocks::*;

`include "awb/provides/unix_comm_device.bsh"

typedef UNIX_COMM_DRIVER SIMULATION_COMMUNICATION_DRIVER;
typedef UNIX_COMM_WIRES  SIMULATION_COMMUNICATION_WIRES;
typedef UNIX_COMM_DEVICE SIMULATION_COMMUNICATION_DEVICE;

module mkSimulationCommunicationDevice#(String outgoing, String incoming) (SIMULATION_COMMUNICATION_DEVICE);
    let commDevice <- mkUNIXCommDevice(outgoing, incoming);
    return commDevice;
endmodule
