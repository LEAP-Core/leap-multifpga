`include "asim/provides/soft_connections.bsh"
`include "asim/provides/test_c.bsh"

module [CONNECTED_MODULE] mkA (Empty);
  let c <- mkC();
endmodule

